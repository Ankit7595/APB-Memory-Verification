class apb_sqr extends uvm_sequencer#(apb_tx);
  
  
  `uvm_component_utils(apb_sqr)
  
      function new (string name="",uvm_component parent=null);
        super.new(name,parent);
      endfunction
      
      function void build_phase (uvm_phase phase);
        super.build_phase(phase);
        $display("apb_sqr::build_phase");
      endfunction 
 endclass